`ifndef PRIM_ASSERT_SV
`define PRIM_ASSERT_SV

`define ASSERT_IF(a1, a2, a3)
`define ASSERT(a1, a2)
`define ASSERT_KNOWN(a1, a2)
`define ASSERT_KNOWN_IF(a1, a2, a3)
`define ASSERT_INIT(a1, a2)

`endif // PRIM_ASSERT_SV
