`ifndef DV_FCOV_MACROS_SVH
`define DV_FCOV_MACROS_SVH

`define DV_FCOV_SIGNAL(a1, a2, a3)
`define DV_FCOV_SIGNAL_GEN_IF(a1, a2, a3, a4)

`endif // DV_FCOV_MACROS_SVH
